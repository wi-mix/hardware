-- soc_system.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		adc_external_interface_sclk         : out   std_logic;                                        --       adc_external_interface.sclk
		adc_external_interface_cs_n         : out   std_logic;                                        --                             .cs_n
		adc_external_interface_dout         : in    std_logic                     := '0';             --                             .dout
		adc_external_interface_din          : out   std_logic;                                        --                             .din
		clk_clk                             : in    std_logic                     := '0';             --                          clk.clk
		hex0_export                         : out   std_logic_vector(6 downto 0);                     --                         hex0.export
		hex1_export                         : out   std_logic_vector(6 downto 0);                     --                         hex1.export
		hex2_export                         : out   std_logic_vector(6 downto 0);                     --                         hex2.export
		hex3_export                         : out   std_logic_vector(6 downto 0);                     --                         hex3.export
		hex4_export                         : out   std_logic_vector(6 downto 0);                     --                         hex4.export
		hex5_export                         : out   std_logic_vector(6 downto 0);                     --                         hex5.export
		hps_io_hps_io_emac1_inst_TX_CLK     : out   std_logic;                                        --                       hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0       : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1       : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2       : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3       : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0       : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO       : inout std_logic                     := '0';             --                             .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC        : out   std_logic;                                        --                             .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL     : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL     : out   std_logic;                                        --                             .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK     : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1       : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2       : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3       : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD3
		hps_io_hps_io_sdio_inst_CMD         : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0          : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1          : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK         : out   std_logic;                                        --                             .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2          : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3          : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7          : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK         : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP         : out   std_logic;                                        --                             .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR         : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT         : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim1_inst_CLK        : out   std_logic;                                        --                             .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI       : out   std_logic;                                        --                             .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO       : in    std_logic                     := '0';             --                             .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0        : out   std_logic;                                        --                             .hps_io_spim1_inst_SS0
		hps_io_hps_io_uart0_inst_RX         : in    std_logic                     := '0';             --                             .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX         : out   std_logic;                                        --                             .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA         : inout std_logic                     := '0';             --                             .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL         : inout std_logic                     := '0';             --                             .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA         : inout std_logic                     := '0';             --                             .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL         : inout std_logic                     := '0';             --                             .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO40      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO48      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO53
		hps_io_hps_io_gpio_inst_GPIO54      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO54
		hps_io_hps_io_gpio_inst_GPIO61      : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO61
		memory_mem_a                        : out   std_logic_vector(14 downto 0);                    --                       memory.mem_a
		memory_mem_ba                       : out   std_logic_vector(2 downto 0);                     --                             .mem_ba
		memory_mem_ck                       : out   std_logic;                                        --                             .mem_ck
		memory_mem_ck_n                     : out   std_logic;                                        --                             .mem_ck_n
		memory_mem_cke                      : out   std_logic;                                        --                             .mem_cke
		memory_mem_cs_n                     : out   std_logic;                                        --                             .mem_cs_n
		memory_mem_ras_n                    : out   std_logic;                                        --                             .mem_ras_n
		memory_mem_cas_n                    : out   std_logic;                                        --                             .mem_cas_n
		memory_mem_we_n                     : out   std_logic;                                        --                             .mem_we_n
		memory_mem_reset_n                  : out   std_logic;                                        --                             .mem_reset_n
		memory_mem_dq                       : inout std_logic_vector(31 downto 0) := (others => '0'); --                             .mem_dq
		memory_mem_dqs                      : inout std_logic_vector(3 downto 0)  := (others => '0'); --                             .mem_dqs
		memory_mem_dqs_n                    : inout std_logic_vector(3 downto 0)  := (others => '0'); --                             .mem_dqs_n
		memory_mem_odt                      : out   std_logic;                                        --                             .mem_odt
		memory_mem_dm                       : out   std_logic_vector(3 downto 0);                     --                             .mem_dm
		memory_oct_rzqin                    : in    std_logic                     := '0';             --                             .oct_rzqin
		multi_pwm_export_pwm1               : out   std_logic;                                        --                    multi_pwm.export_pwm1
		multi_pwm_export_pwm2               : out   std_logic;                                        --                             .export_pwm2
		multi_pwm_export_pwm3               : out   std_logic;                                        --                             .export_pwm3
		multi_pwm_export_pwm4               : out   std_logic;                                        --                             .export_pwm4
		red_leds_external_connection_export : out   std_logic_vector(9 downto 0);                     -- red_leds_external_connection.export
		reset_reset_n                       : in    std_logic                     := '0';             --                        reset.reset_n
		switches_external_connection_export : in    std_logic_vector(9 downto 0)  := (others => '0')  -- switches_external_connection.export
	);
end entity soc_system;

architecture rtl of soc_system is
	component soc_system_adc is
		generic (
			board          : string  := "DE10-Standard";
			board_rev      : string  := "Autodetect";
			tsclk          : integer := 0;
			numch          : integer := 0;
			max10pllmultby : integer := 0;
			max10plldivby  : integer := 0
		);
		port (
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			waitrequest : out std_logic;                                        -- waitrequest
			read        : in  std_logic                     := 'X';             -- read
			adc_sclk    : out std_logic;                                        -- export
			adc_cs_n    : out std_logic;                                        -- export
			adc_dout    : in  std_logic                     := 'X';             -- export
			adc_din     : out std_logic                                         -- export
		);
	end component soc_system_adc;

	component seven_seg is
		port (
			avalon_slave_write_n   : in  std_logic                     := 'X';             -- write_n
			avalon_slave_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clk                    : in  std_logic                     := 'X';             -- clk
			conduit_end_hex        : out std_logic_vector(6 downto 0);                     -- export
			reset_n                : in  std_logic                     := 'X'              -- reset_n
		);
	end component seven_seg;

	component soc_system_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                         -- rready
		);
	end component soc_system_hps;

	component multi_pwm is
		generic (
			W : integer := 15
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset_n   : in  std_logic                     := 'X';             -- reset_n
			writas    : in  std_logic                     := 'X';             -- write_n
			address   : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			PWM1      : out std_logic;                                        -- export_pwm1
			PWM2      : out std_logic;                                        -- export_pwm2
			PWM3      : out std_logic;                                        -- export_pwm3
			PWM4      : out std_logic                                         -- export_pwm4
		);
	end component multi_pwm;

	component soc_system_red_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component soc_system_red_leds;

	component soc_system_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component soc_system_switches;

	component soc_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid_qsys_0;

	component soc_system_mm_interconnect_0 is
		port (
			hps_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                     : in  std_logic                     := 'X';             -- clk
			adc_reset_reset_bridge_in_reset_reset                             : in  std_logic                     := 'X';             -- reset
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			adc_adc_slave_address                                             : out std_logic_vector(2 downto 0);                     -- address
			adc_adc_slave_write                                               : out std_logic;                                        -- write
			adc_adc_slave_read                                                : out std_logic;                                        -- read
			adc_adc_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			adc_adc_slave_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			adc_adc_slave_waitrequest                                         : in  std_logic                     := 'X';             -- waitrequest
			hex0_avalon_slave_write                                           : out std_logic;                                        -- write
			hex0_avalon_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex1_avalon_slave_write                                           : out std_logic;                                        -- write
			hex1_avalon_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex2_avalon_slave_write                                           : out std_logic;                                        -- write
			hex2_avalon_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex3_avalon_slave_write                                           : out std_logic;                                        -- write
			hex3_avalon_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex4_avalon_slave_write                                           : out std_logic;                                        -- write
			hex4_avalon_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			hex5_avalon_slave_write                                           : out std_logic;                                        -- write
			hex5_avalon_slave_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			multi_pwm_0_avalon_slave_0_address                                : out std_logic_vector(5 downto 0);                     -- address
			multi_pwm_0_avalon_slave_0_write                                  : out std_logic;                                        -- write
			multi_pwm_0_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			red_leds_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			red_leds_s1_write                                                 : out std_logic;                                        -- write
			red_leds_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			red_leds_s1_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			red_leds_s1_chipselect                                            : out std_logic;                                        -- chipselect
			switches_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_0_control_slave_address                                : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	signal hps_h2f_lw_axi_master_awburst                                : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_awburst
	signal hps_h2f_lw_axi_master_arlen                                  : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_arlen
	signal hps_h2f_lw_axi_master_wstrb                                  : std_logic_vector(3 downto 0);  -- hps:h2f_lw_WSTRB -> mm_interconnect_0:hps_h2f_lw_axi_master_wstrb
	signal hps_h2f_lw_axi_master_wready                                 : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	signal hps_h2f_lw_axi_master_rid                                    : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	signal hps_h2f_lw_axi_master_rready                                 : std_logic;                     -- hps:h2f_lw_RREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_rready
	signal hps_h2f_lw_axi_master_awlen                                  : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_awlen
	signal hps_h2f_lw_axi_master_wid                                    : std_logic_vector(11 downto 0); -- hps:h2f_lw_WID -> mm_interconnect_0:hps_h2f_lw_axi_master_wid
	signal hps_h2f_lw_axi_master_arcache                                : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_arcache
	signal hps_h2f_lw_axi_master_wvalid                                 : std_logic;                     -- hps:h2f_lw_WVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_wvalid
	signal hps_h2f_lw_axi_master_araddr                                 : std_logic_vector(20 downto 0); -- hps:h2f_lw_ARADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_araddr
	signal hps_h2f_lw_axi_master_arprot                                 : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_arprot
	signal hps_h2f_lw_axi_master_awprot                                 : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_awprot
	signal hps_h2f_lw_axi_master_wdata                                  : std_logic_vector(31 downto 0); -- hps:h2f_lw_WDATA -> mm_interconnect_0:hps_h2f_lw_axi_master_wdata
	signal hps_h2f_lw_axi_master_arvalid                                : std_logic;                     -- hps:h2f_lw_ARVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_arvalid
	signal hps_h2f_lw_axi_master_awcache                                : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_awcache
	signal hps_h2f_lw_axi_master_arid                                   : std_logic_vector(11 downto 0); -- hps:h2f_lw_ARID -> mm_interconnect_0:hps_h2f_lw_axi_master_arid
	signal hps_h2f_lw_axi_master_arlock                                 : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_arlock
	signal hps_h2f_lw_axi_master_awlock                                 : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_awlock
	signal hps_h2f_lw_axi_master_awaddr                                 : std_logic_vector(20 downto 0); -- hps:h2f_lw_AWADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_awaddr
	signal hps_h2f_lw_axi_master_bresp                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	signal hps_h2f_lw_axi_master_arready                                : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	signal hps_h2f_lw_axi_master_rdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	signal hps_h2f_lw_axi_master_awready                                : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	signal hps_h2f_lw_axi_master_arburst                                : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_arburst
	signal hps_h2f_lw_axi_master_arsize                                 : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_arsize
	signal hps_h2f_lw_axi_master_bready                                 : std_logic;                     -- hps:h2f_lw_BREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_bready
	signal hps_h2f_lw_axi_master_rlast                                  : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	signal hps_h2f_lw_axi_master_wlast                                  : std_logic;                     -- hps:h2f_lw_WLAST -> mm_interconnect_0:hps_h2f_lw_axi_master_wlast
	signal hps_h2f_lw_axi_master_rresp                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	signal hps_h2f_lw_axi_master_awid                                   : std_logic_vector(11 downto 0); -- hps:h2f_lw_AWID -> mm_interconnect_0:hps_h2f_lw_axi_master_awid
	signal hps_h2f_lw_axi_master_bid                                    : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	signal hps_h2f_lw_axi_master_bvalid                                 : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	signal hps_h2f_lw_axi_master_awsize                                 : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_awsize
	signal hps_h2f_lw_axi_master_awvalid                                : std_logic;                     -- hps:h2f_lw_AWVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_awvalid
	signal hps_h2f_lw_axi_master_rvalid                                 : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	signal mm_interconnect_0_adc_adc_slave_readdata                     : std_logic_vector(31 downto 0); -- adc:readdata -> mm_interconnect_0:adc_adc_slave_readdata
	signal mm_interconnect_0_adc_adc_slave_waitrequest                  : std_logic;                     -- adc:waitrequest -> mm_interconnect_0:adc_adc_slave_waitrequest
	signal mm_interconnect_0_adc_adc_slave_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:adc_adc_slave_address -> adc:address
	signal mm_interconnect_0_adc_adc_slave_read                         : std_logic;                     -- mm_interconnect_0:adc_adc_slave_read -> adc:read
	signal mm_interconnect_0_adc_adc_slave_write                        : std_logic;                     -- mm_interconnect_0:adc_adc_slave_write -> adc:write
	signal mm_interconnect_0_adc_adc_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:adc_adc_slave_writedata -> adc:writedata
	signal mm_interconnect_0_hex0_avalon_slave_write                    : std_logic;                     -- mm_interconnect_0:hex0_avalon_slave_write -> mm_interconnect_0_hex0_avalon_slave_write:in
	signal mm_interconnect_0_hex0_avalon_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex0_avalon_slave_writedata -> hex0:avalon_slave_writedata
	signal mm_interconnect_0_hex1_avalon_slave_write                    : std_logic;                     -- mm_interconnect_0:hex1_avalon_slave_write -> mm_interconnect_0_hex1_avalon_slave_write:in
	signal mm_interconnect_0_hex1_avalon_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex1_avalon_slave_writedata -> hex1:avalon_slave_writedata
	signal mm_interconnect_0_hex2_avalon_slave_write                    : std_logic;                     -- mm_interconnect_0:hex2_avalon_slave_write -> mm_interconnect_0_hex2_avalon_slave_write:in
	signal mm_interconnect_0_hex2_avalon_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex2_avalon_slave_writedata -> hex2:avalon_slave_writedata
	signal mm_interconnect_0_hex3_avalon_slave_write                    : std_logic;                     -- mm_interconnect_0:hex3_avalon_slave_write -> mm_interconnect_0_hex3_avalon_slave_write:in
	signal mm_interconnect_0_hex3_avalon_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex3_avalon_slave_writedata -> hex3:avalon_slave_writedata
	signal mm_interconnect_0_hex4_avalon_slave_write                    : std_logic;                     -- mm_interconnect_0:hex4_avalon_slave_write -> mm_interconnect_0_hex4_avalon_slave_write:in
	signal mm_interconnect_0_hex4_avalon_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex4_avalon_slave_writedata -> hex4:avalon_slave_writedata
	signal mm_interconnect_0_hex5_avalon_slave_write                    : std_logic;                     -- mm_interconnect_0:hex5_avalon_slave_write -> mm_interconnect_0_hex5_avalon_slave_write:in
	signal mm_interconnect_0_hex5_avalon_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex5_avalon_slave_writedata -> hex5:avalon_slave_writedata
	signal mm_interconnect_0_multi_pwm_0_avalon_slave_0_address         : std_logic_vector(5 downto 0);  -- mm_interconnect_0:multi_pwm_0_avalon_slave_0_address -> multi_pwm_0:address
	signal mm_interconnect_0_multi_pwm_0_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:multi_pwm_0_avalon_slave_0_write -> mm_interconnect_0_multi_pwm_0_avalon_slave_0_write:in
	signal mm_interconnect_0_multi_pwm_0_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:multi_pwm_0_avalon_slave_0_writedata -> multi_pwm_0:writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata        : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_red_leds_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:red_leds_s1_chipselect -> red_leds:chipselect
	signal mm_interconnect_0_red_leds_s1_readdata                       : std_logic_vector(31 downto 0); -- red_leds:readdata -> mm_interconnect_0:red_leds_s1_readdata
	signal mm_interconnect_0_red_leds_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:red_leds_s1_address -> red_leds:address
	signal mm_interconnect_0_red_leds_s1_write                          : std_logic;                     -- mm_interconnect_0:red_leds_s1_write -> mm_interconnect_0_red_leds_s1_write:in
	signal mm_interconnect_0_red_leds_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_leds_s1_writedata -> red_leds:writedata
	signal mm_interconnect_0_switches_s1_readdata                       : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [adc:reset, mm_interconnect_0:adc_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal hps_h2f_reset_reset                                          : std_logic;                     -- hps:h2f_rst_n -> hps_h2f_reset_reset:in
	signal rst_controller_001_reset_out_reset                           : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_0:hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal reset_reset_n_ports_inv                                      : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_hex0_avalon_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_hex0_avalon_slave_write:inv -> hex0:avalon_slave_write_n
	signal mm_interconnect_0_hex1_avalon_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_hex1_avalon_slave_write:inv -> hex1:avalon_slave_write_n
	signal mm_interconnect_0_hex2_avalon_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_hex2_avalon_slave_write:inv -> hex2:avalon_slave_write_n
	signal mm_interconnect_0_hex3_avalon_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_hex3_avalon_slave_write:inv -> hex3:avalon_slave_write_n
	signal mm_interconnect_0_hex4_avalon_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_hex4_avalon_slave_write:inv -> hex4:avalon_slave_write_n
	signal mm_interconnect_0_hex5_avalon_slave_write_ports_inv          : std_logic;                     -- mm_interconnect_0_hex5_avalon_slave_write:inv -> hex5:avalon_slave_write_n
	signal mm_interconnect_0_multi_pwm_0_avalon_slave_0_write_ports_inv : std_logic;                     -- mm_interconnect_0_multi_pwm_0_avalon_slave_0_write:inv -> multi_pwm_0:writas
	signal mm_interconnect_0_red_leds_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_red_leds_s1_write:inv -> red_leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> [hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, multi_pwm_0:reset_n, red_leds:reset_n, switches:reset_n, sysid_qsys_0:reset_n]
	signal hps_h2f_reset_reset_ports_inv                                : std_logic;                     -- hps_h2f_reset_reset:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in0]

begin

	adc : component soc_system_adc
		generic map (
			board          => "DE1-SoC",
			board_rev      => "F or newer",
			tsclk          => 4,
			numch          => 7,
			max10pllmultby => 1,
			max10plldivby  => 1
		)
		port map (
			clock       => clk_clk,                                     --                clk.clk
			reset       => rst_controller_reset_out_reset,              --              reset.reset
			write       => mm_interconnect_0_adc_adc_slave_write,       --          adc_slave.write
			readdata    => mm_interconnect_0_adc_adc_slave_readdata,    --                   .readdata
			writedata   => mm_interconnect_0_adc_adc_slave_writedata,   --                   .writedata
			address     => mm_interconnect_0_adc_adc_slave_address,     --                   .address
			waitrequest => mm_interconnect_0_adc_adc_slave_waitrequest, --                   .waitrequest
			read        => mm_interconnect_0_adc_adc_slave_read,        --                   .read
			adc_sclk    => adc_external_interface_sclk,                 -- external_interface.export
			adc_cs_n    => adc_external_interface_cs_n,                 --                   .export
			adc_dout    => adc_external_interface_dout,                 --                   .export
			adc_din     => adc_external_interface_din                   --                   .export
		);

	hex0 : component seven_seg
		port map (
			avalon_slave_write_n   => mm_interconnect_0_hex0_avalon_slave_write_ports_inv, -- avalon_slave.write_n
			avalon_slave_writedata => mm_interconnect_0_hex0_avalon_slave_writedata,       --             .writedata
			clk                    => clk_clk,                                             --        clock.clk
			conduit_end_hex        => hex0_export,                                         --      conduit.export
			reset_n                => rst_controller_reset_out_reset_ports_inv             --        reset.reset_n
		);

	hex1 : component seven_seg
		port map (
			avalon_slave_write_n   => mm_interconnect_0_hex1_avalon_slave_write_ports_inv, -- avalon_slave.write_n
			avalon_slave_writedata => mm_interconnect_0_hex1_avalon_slave_writedata,       --             .writedata
			clk                    => clk_clk,                                             --        clock.clk
			conduit_end_hex        => hex1_export,                                         --      conduit.export
			reset_n                => rst_controller_reset_out_reset_ports_inv             --        reset.reset_n
		);

	hex2 : component seven_seg
		port map (
			avalon_slave_write_n   => mm_interconnect_0_hex2_avalon_slave_write_ports_inv, -- avalon_slave.write_n
			avalon_slave_writedata => mm_interconnect_0_hex2_avalon_slave_writedata,       --             .writedata
			clk                    => clk_clk,                                             --        clock.clk
			conduit_end_hex        => hex2_export,                                         --      conduit.export
			reset_n                => rst_controller_reset_out_reset_ports_inv             --        reset.reset_n
		);

	hex3 : component seven_seg
		port map (
			avalon_slave_write_n   => mm_interconnect_0_hex3_avalon_slave_write_ports_inv, -- avalon_slave.write_n
			avalon_slave_writedata => mm_interconnect_0_hex3_avalon_slave_writedata,       --             .writedata
			clk                    => clk_clk,                                             --        clock.clk
			conduit_end_hex        => hex3_export,                                         --      conduit.export
			reset_n                => rst_controller_reset_out_reset_ports_inv             --        reset.reset_n
		);

	hex4 : component seven_seg
		port map (
			avalon_slave_write_n   => mm_interconnect_0_hex4_avalon_slave_write_ports_inv, -- avalon_slave.write_n
			avalon_slave_writedata => mm_interconnect_0_hex4_avalon_slave_writedata,       --             .writedata
			clk                    => clk_clk,                                             --        clock.clk
			conduit_end_hex        => hex4_export,                                         --      conduit.export
			reset_n                => rst_controller_reset_out_reset_ports_inv             --        reset.reset_n
		);

	hex5 : component seven_seg
		port map (
			avalon_slave_write_n   => mm_interconnect_0_hex5_avalon_slave_write_ports_inv, -- avalon_slave.write_n
			avalon_slave_writedata => mm_interconnect_0_hex5_avalon_slave_writedata,       --             .writedata
			clk                    => clk_clk,                                             --        clock.clk
			conduit_end_hex        => hex5_export,                                         --      conduit.export
			reset_n                => rst_controller_reset_out_reset_ports_inv             --        reset.reset_n
		);

	hps : component soc_system_hps
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => memory_mem_a,                    --            memory.mem_a
			mem_ba                   => memory_mem_ba,                   --                  .mem_ba
			mem_ck                   => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                  --                  .mem_odt
			mem_dm                   => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK, --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,   --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,   --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,   --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,   --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,   --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,   --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,    --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL, --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL, --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK, --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,   --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,   --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,   --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,     --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,      --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,      --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,     --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,      --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,      --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,      --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,      --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,      --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,      --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,      --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,      --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,      --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,      --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,     --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,     --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,     --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,     --                  .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_io_hps_io_spim1_inst_CLK,    --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_io_hps_io_spim1_inst_MOSI,   --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_io_hps_io_spim1_inst_MISO,   --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_io_hps_io_spim1_inst_SS0,    --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,     --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,     --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,     --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,     --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,     --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_io_hps_io_gpio_inst_GPIO09,  --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_io_hps_io_gpio_inst_GPIO35,  --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_io_hps_io_gpio_inst_GPIO40,  --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  => hps_io_hps_io_gpio_inst_GPIO48,  --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_io_hps_io_gpio_inst_GPIO53,  --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_io_hps_io_gpio_inst_GPIO54,  --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_io_hps_io_gpio_inst_GPIO61,  --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_h2f_reset_reset,             --         h2f_reset.reset_n
			h2f_lw_axi_clk           => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_h2f_lw_axi_master_awid,      -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_h2f_lw_axi_master_awaddr,    --                  .awaddr
			h2f_lw_AWLEN             => hps_h2f_lw_axi_master_awlen,     --                  .awlen
			h2f_lw_AWSIZE            => hps_h2f_lw_axi_master_awsize,    --                  .awsize
			h2f_lw_AWBURST           => hps_h2f_lw_axi_master_awburst,   --                  .awburst
			h2f_lw_AWLOCK            => hps_h2f_lw_axi_master_awlock,    --                  .awlock
			h2f_lw_AWCACHE           => hps_h2f_lw_axi_master_awcache,   --                  .awcache
			h2f_lw_AWPROT            => hps_h2f_lw_axi_master_awprot,    --                  .awprot
			h2f_lw_AWVALID           => hps_h2f_lw_axi_master_awvalid,   --                  .awvalid
			h2f_lw_AWREADY           => hps_h2f_lw_axi_master_awready,   --                  .awready
			h2f_lw_WID               => hps_h2f_lw_axi_master_wid,       --                  .wid
			h2f_lw_WDATA             => hps_h2f_lw_axi_master_wdata,     --                  .wdata
			h2f_lw_WSTRB             => hps_h2f_lw_axi_master_wstrb,     --                  .wstrb
			h2f_lw_WLAST             => hps_h2f_lw_axi_master_wlast,     --                  .wlast
			h2f_lw_WVALID            => hps_h2f_lw_axi_master_wvalid,    --                  .wvalid
			h2f_lw_WREADY            => hps_h2f_lw_axi_master_wready,    --                  .wready
			h2f_lw_BID               => hps_h2f_lw_axi_master_bid,       --                  .bid
			h2f_lw_BRESP             => hps_h2f_lw_axi_master_bresp,     --                  .bresp
			h2f_lw_BVALID            => hps_h2f_lw_axi_master_bvalid,    --                  .bvalid
			h2f_lw_BREADY            => hps_h2f_lw_axi_master_bready,    --                  .bready
			h2f_lw_ARID              => hps_h2f_lw_axi_master_arid,      --                  .arid
			h2f_lw_ARADDR            => hps_h2f_lw_axi_master_araddr,    --                  .araddr
			h2f_lw_ARLEN             => hps_h2f_lw_axi_master_arlen,     --                  .arlen
			h2f_lw_ARSIZE            => hps_h2f_lw_axi_master_arsize,    --                  .arsize
			h2f_lw_ARBURST           => hps_h2f_lw_axi_master_arburst,   --                  .arburst
			h2f_lw_ARLOCK            => hps_h2f_lw_axi_master_arlock,    --                  .arlock
			h2f_lw_ARCACHE           => hps_h2f_lw_axi_master_arcache,   --                  .arcache
			h2f_lw_ARPROT            => hps_h2f_lw_axi_master_arprot,    --                  .arprot
			h2f_lw_ARVALID           => hps_h2f_lw_axi_master_arvalid,   --                  .arvalid
			h2f_lw_ARREADY           => hps_h2f_lw_axi_master_arready,   --                  .arready
			h2f_lw_RID               => hps_h2f_lw_axi_master_rid,       --                  .rid
			h2f_lw_RDATA             => hps_h2f_lw_axi_master_rdata,     --                  .rdata
			h2f_lw_RRESP             => hps_h2f_lw_axi_master_rresp,     --                  .rresp
			h2f_lw_RLAST             => hps_h2f_lw_axi_master_rlast,     --                  .rlast
			h2f_lw_RVALID            => hps_h2f_lw_axi_master_rvalid,    --                  .rvalid
			h2f_lw_RREADY            => hps_h2f_lw_axi_master_rready     --                  .rready
		);

	multi_pwm_0 : component multi_pwm
		generic map (
			W => 31
		)
		port map (
			clk       => clk_clk,                                                      --          clock.clk
			reset_n   => rst_controller_reset_out_reset_ports_inv,                     --          reset.reset_n
			writas    => mm_interconnect_0_multi_pwm_0_avalon_slave_0_write_ports_inv, -- avalon_slave_0.write_n
			address   => mm_interconnect_0_multi_pwm_0_avalon_slave_0_address,         --               .address
			writedata => mm_interconnect_0_multi_pwm_0_avalon_slave_0_writedata,       --               .writedata
			PWM1      => multi_pwm_export_pwm1,                                        --    conduit_end.export_pwm1
			PWM2      => multi_pwm_export_pwm2,                                        --               .export_pwm2
			PWM3      => multi_pwm_export_pwm3,                                        --               .export_pwm3
			PWM4      => multi_pwm_export_pwm4                                         --               .export_pwm4
		);

	red_leds : component soc_system_red_leds
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_red_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_red_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_red_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_red_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_red_leds_s1_readdata,        --                    .readdata
			out_port   => red_leds_external_connection_export            -- external_connection.export
		);

	switches : component soc_system_switches
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,   --                    .readdata
			in_port  => switches_external_connection_export       -- external_connection.export
		);

	sysid_qsys_0 : component soc_system_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			hps_h2f_lw_axi_master_awid                                        => hps_h2f_lw_axi_master_awid,                             --                                       hps_h2f_lw_axi_master.awid
			hps_h2f_lw_axi_master_awaddr                                      => hps_h2f_lw_axi_master_awaddr,                           --                                                            .awaddr
			hps_h2f_lw_axi_master_awlen                                       => hps_h2f_lw_axi_master_awlen,                            --                                                            .awlen
			hps_h2f_lw_axi_master_awsize                                      => hps_h2f_lw_axi_master_awsize,                           --                                                            .awsize
			hps_h2f_lw_axi_master_awburst                                     => hps_h2f_lw_axi_master_awburst,                          --                                                            .awburst
			hps_h2f_lw_axi_master_awlock                                      => hps_h2f_lw_axi_master_awlock,                           --                                                            .awlock
			hps_h2f_lw_axi_master_awcache                                     => hps_h2f_lw_axi_master_awcache,                          --                                                            .awcache
			hps_h2f_lw_axi_master_awprot                                      => hps_h2f_lw_axi_master_awprot,                           --                                                            .awprot
			hps_h2f_lw_axi_master_awvalid                                     => hps_h2f_lw_axi_master_awvalid,                          --                                                            .awvalid
			hps_h2f_lw_axi_master_awready                                     => hps_h2f_lw_axi_master_awready,                          --                                                            .awready
			hps_h2f_lw_axi_master_wid                                         => hps_h2f_lw_axi_master_wid,                              --                                                            .wid
			hps_h2f_lw_axi_master_wdata                                       => hps_h2f_lw_axi_master_wdata,                            --                                                            .wdata
			hps_h2f_lw_axi_master_wstrb                                       => hps_h2f_lw_axi_master_wstrb,                            --                                                            .wstrb
			hps_h2f_lw_axi_master_wlast                                       => hps_h2f_lw_axi_master_wlast,                            --                                                            .wlast
			hps_h2f_lw_axi_master_wvalid                                      => hps_h2f_lw_axi_master_wvalid,                           --                                                            .wvalid
			hps_h2f_lw_axi_master_wready                                      => hps_h2f_lw_axi_master_wready,                           --                                                            .wready
			hps_h2f_lw_axi_master_bid                                         => hps_h2f_lw_axi_master_bid,                              --                                                            .bid
			hps_h2f_lw_axi_master_bresp                                       => hps_h2f_lw_axi_master_bresp,                            --                                                            .bresp
			hps_h2f_lw_axi_master_bvalid                                      => hps_h2f_lw_axi_master_bvalid,                           --                                                            .bvalid
			hps_h2f_lw_axi_master_bready                                      => hps_h2f_lw_axi_master_bready,                           --                                                            .bready
			hps_h2f_lw_axi_master_arid                                        => hps_h2f_lw_axi_master_arid,                             --                                                            .arid
			hps_h2f_lw_axi_master_araddr                                      => hps_h2f_lw_axi_master_araddr,                           --                                                            .araddr
			hps_h2f_lw_axi_master_arlen                                       => hps_h2f_lw_axi_master_arlen,                            --                                                            .arlen
			hps_h2f_lw_axi_master_arsize                                      => hps_h2f_lw_axi_master_arsize,                           --                                                            .arsize
			hps_h2f_lw_axi_master_arburst                                     => hps_h2f_lw_axi_master_arburst,                          --                                                            .arburst
			hps_h2f_lw_axi_master_arlock                                      => hps_h2f_lw_axi_master_arlock,                           --                                                            .arlock
			hps_h2f_lw_axi_master_arcache                                     => hps_h2f_lw_axi_master_arcache,                          --                                                            .arcache
			hps_h2f_lw_axi_master_arprot                                      => hps_h2f_lw_axi_master_arprot,                           --                                                            .arprot
			hps_h2f_lw_axi_master_arvalid                                     => hps_h2f_lw_axi_master_arvalid,                          --                                                            .arvalid
			hps_h2f_lw_axi_master_arready                                     => hps_h2f_lw_axi_master_arready,                          --                                                            .arready
			hps_h2f_lw_axi_master_rid                                         => hps_h2f_lw_axi_master_rid,                              --                                                            .rid
			hps_h2f_lw_axi_master_rdata                                       => hps_h2f_lw_axi_master_rdata,                            --                                                            .rdata
			hps_h2f_lw_axi_master_rresp                                       => hps_h2f_lw_axi_master_rresp,                            --                                                            .rresp
			hps_h2f_lw_axi_master_rlast                                       => hps_h2f_lw_axi_master_rlast,                            --                                                            .rlast
			hps_h2f_lw_axi_master_rvalid                                      => hps_h2f_lw_axi_master_rvalid,                           --                                                            .rvalid
			hps_h2f_lw_axi_master_rready                                      => hps_h2f_lw_axi_master_rready,                           --                                                            .rready
			clk_0_clk_clk                                                     => clk_clk,                                                --                                                   clk_0_clk.clk
			adc_reset_reset_bridge_in_reset_reset                             => rst_controller_reset_out_reset,                         --                             adc_reset_reset_bridge_in_reset.reset
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                     -- hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			adc_adc_slave_address                                             => mm_interconnect_0_adc_adc_slave_address,                --                                               adc_adc_slave.address
			adc_adc_slave_write                                               => mm_interconnect_0_adc_adc_slave_write,                  --                                                            .write
			adc_adc_slave_read                                                => mm_interconnect_0_adc_adc_slave_read,                   --                                                            .read
			adc_adc_slave_readdata                                            => mm_interconnect_0_adc_adc_slave_readdata,               --                                                            .readdata
			adc_adc_slave_writedata                                           => mm_interconnect_0_adc_adc_slave_writedata,              --                                                            .writedata
			adc_adc_slave_waitrequest                                         => mm_interconnect_0_adc_adc_slave_waitrequest,            --                                                            .waitrequest
			hex0_avalon_slave_write                                           => mm_interconnect_0_hex0_avalon_slave_write,              --                                           hex0_avalon_slave.write
			hex0_avalon_slave_writedata                                       => mm_interconnect_0_hex0_avalon_slave_writedata,          --                                                            .writedata
			hex1_avalon_slave_write                                           => mm_interconnect_0_hex1_avalon_slave_write,              --                                           hex1_avalon_slave.write
			hex1_avalon_slave_writedata                                       => mm_interconnect_0_hex1_avalon_slave_writedata,          --                                                            .writedata
			hex2_avalon_slave_write                                           => mm_interconnect_0_hex2_avalon_slave_write,              --                                           hex2_avalon_slave.write
			hex2_avalon_slave_writedata                                       => mm_interconnect_0_hex2_avalon_slave_writedata,          --                                                            .writedata
			hex3_avalon_slave_write                                           => mm_interconnect_0_hex3_avalon_slave_write,              --                                           hex3_avalon_slave.write
			hex3_avalon_slave_writedata                                       => mm_interconnect_0_hex3_avalon_slave_writedata,          --                                                            .writedata
			hex4_avalon_slave_write                                           => mm_interconnect_0_hex4_avalon_slave_write,              --                                           hex4_avalon_slave.write
			hex4_avalon_slave_writedata                                       => mm_interconnect_0_hex4_avalon_slave_writedata,          --                                                            .writedata
			hex5_avalon_slave_write                                           => mm_interconnect_0_hex5_avalon_slave_write,              --                                           hex5_avalon_slave.write
			hex5_avalon_slave_writedata                                       => mm_interconnect_0_hex5_avalon_slave_writedata,          --                                                            .writedata
			multi_pwm_0_avalon_slave_0_address                                => mm_interconnect_0_multi_pwm_0_avalon_slave_0_address,   --                                  multi_pwm_0_avalon_slave_0.address
			multi_pwm_0_avalon_slave_0_write                                  => mm_interconnect_0_multi_pwm_0_avalon_slave_0_write,     --                                                            .write
			multi_pwm_0_avalon_slave_0_writedata                              => mm_interconnect_0_multi_pwm_0_avalon_slave_0_writedata, --                                                            .writedata
			red_leds_s1_address                                               => mm_interconnect_0_red_leds_s1_address,                  --                                                 red_leds_s1.address
			red_leds_s1_write                                                 => mm_interconnect_0_red_leds_s1_write,                    --                                                            .write
			red_leds_s1_readdata                                              => mm_interconnect_0_red_leds_s1_readdata,                 --                                                            .readdata
			red_leds_s1_writedata                                             => mm_interconnect_0_red_leds_s1_writedata,                --                                                            .writedata
			red_leds_s1_chipselect                                            => mm_interconnect_0_red_leds_s1_chipselect,               --                                                            .chipselect
			switches_s1_address                                               => mm_interconnect_0_switches_s1_address,                  --                                                 switches_s1.address
			switches_s1_readdata                                              => mm_interconnect_0_switches_s1_readdata,                 --                                                            .readdata
			sysid_qsys_0_control_slave_address                                => mm_interconnect_0_sysid_qsys_0_control_slave_address,   --                                  sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                               => mm_interconnect_0_sysid_qsys_0_control_slave_readdata   --                                                            .readdata
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			reset_in1      => hps_h2f_reset_reset_ports_inv,  -- reset_in1.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_h2f_reset_reset_ports_inv,      -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_hex0_avalon_slave_write_ports_inv <= not mm_interconnect_0_hex0_avalon_slave_write;

	mm_interconnect_0_hex1_avalon_slave_write_ports_inv <= not mm_interconnect_0_hex1_avalon_slave_write;

	mm_interconnect_0_hex2_avalon_slave_write_ports_inv <= not mm_interconnect_0_hex2_avalon_slave_write;

	mm_interconnect_0_hex3_avalon_slave_write_ports_inv <= not mm_interconnect_0_hex3_avalon_slave_write;

	mm_interconnect_0_hex4_avalon_slave_write_ports_inv <= not mm_interconnect_0_hex4_avalon_slave_write;

	mm_interconnect_0_hex5_avalon_slave_write_ports_inv <= not mm_interconnect_0_hex5_avalon_slave_write;

	mm_interconnect_0_multi_pwm_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_multi_pwm_0_avalon_slave_0_write;

	mm_interconnect_0_red_leds_s1_write_ports_inv <= not mm_interconnect_0_red_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_h2f_reset_reset_ports_inv <= not hps_h2f_reset_reset;

end architecture rtl; -- of soc_system
